`include "spi_defines.svh" // For macros
import shared_pkg::*; // For enums and parameters

module golden_model (
    input logic clk
    );

endmodule
