/*  
    This assertion file follows the **Verification Plan** numbering  
    Each section corresponds to a specific verification requirement

    The numbers (e.g., 1, 2.2) match the corresponding test items  
    from the **Verification Plan** for traceability and clarity
*/
`include "spi_defines.svh" // For macros
import shared_pkg::*; // For enums and parameters
`timescale `TIME_UNIT / `TIME_PRECISION

module SPI_slave_sva(
   
	// input [9:0] din,
	// input clk,rst_n,rx_valid,

	// output logic [ADDR_SIZE-1:0] dout,
	// output logic tx_valid

    );
    
   
endmodule